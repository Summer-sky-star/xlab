// soc_system_top_0.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system_top_0 (
		output wire [31:0]  avmm_1_rw_address,       // avmm_1_rw.address
		output wire [15:0]  avmm_1_rw_byteenable,    //          .byteenable
		input  wire         avmm_1_rw_readdatavalid, //          .readdatavalid
		output wire         avmm_1_rw_read,          //          .read
		input  wire [127:0] avmm_1_rw_readdata,      //          .readdata
		output wire         avmm_1_rw_write,         //          .write
		output wire [127:0] avmm_1_rw_writedata,     //          .writedata
		input  wire         avmm_1_rw_waitrequest,   //          .waitrequest
		output wire         avmm_1_rw_burstcount,    //          .burstcount
		output wire [31:0]  avmm_2_rw_address,       // avmm_2_rw.address
		output wire [15:0]  avmm_2_rw_byteenable,    //          .byteenable
		input  wire         avmm_2_rw_readdatavalid, //          .readdatavalid
		output wire         avmm_2_rw_read,          //          .read
		input  wire [127:0] avmm_2_rw_readdata,      //          .readdata
		output wire         avmm_2_rw_write,         //          .write
		output wire [127:0] avmm_2_rw_writedata,     //          .writedata
		input  wire         avmm_2_rw_waitrequest,   //          .waitrequest
		output wire         avmm_2_rw_burstcount,    //          .burstcount
		output wire [31:0]  avmm_3_rw_address,       // avmm_3_rw.address
		output wire [3:0]   avmm_3_rw_byteenable,    //          .byteenable
		input  wire         avmm_3_rw_readdatavalid, //          .readdatavalid
		output wire         avmm_3_rw_read,          //          .read
		input  wire [31:0]  avmm_3_rw_readdata,      //          .readdata
		output wire         avmm_3_rw_write,         //          .write
		output wire [31:0]  avmm_3_rw_writedata,     //          .writedata
		input  wire         avmm_3_rw_waitrequest,   //          .waitrequest
		output wire         avmm_3_rw_burstcount,    //          .burstcount
		output wire [31:0]  avmm_4_rw_address,       // avmm_4_rw.address
		output wire [3:0]   avmm_4_rw_byteenable,    //          .byteenable
		input  wire         avmm_4_rw_readdatavalid, //          .readdatavalid
		output wire         avmm_4_rw_read,          //          .read
		input  wire [31:0]  avmm_4_rw_readdata,      //          .readdata
		output wire         avmm_4_rw_write,         //          .write
		output wire [31:0]  avmm_4_rw_writedata,     //          .writedata
		input  wire         avmm_4_rw_waitrequest,   //          .waitrequest
		output wire         avmm_4_rw_burstcount,    //          .burstcount
		output wire [31:0]  avmm_5_rw_address,       // avmm_5_rw.address
		output wire [3:0]   avmm_5_rw_byteenable,    //          .byteenable
		input  wire         avmm_5_rw_readdatavalid, //          .readdatavalid
		output wire         avmm_5_rw_read,          //          .read
		input  wire [31:0]  avmm_5_rw_readdata,      //          .readdata
		output wire         avmm_5_rw_write,         //          .write
		output wire [31:0]  avmm_5_rw_writedata,     //          .writedata
		input  wire         avmm_5_rw_waitrequest,   //          .waitrequest
		output wire         avmm_5_rw_burstcount,    //          .burstcount
		input  wire         start,                   //      call.valid
		output wire         busy,                    //          .stall
		input  wire         clock,                   //     clock.clk
		input  wire [63:0]  ddr_in1,                 //   ddr_in1.data
		input  wire [63:0]  ddr_out1,                //  ddr_out1.data
		input  wire [63:0]  ddr_scale,               // ddr_scale.data
		input  wire [63:0]  ddr_w1,                  //    ddr_w1.data
		input  wire [63:0]  param,                   //     param.data
		input  wire         resetn,                  //     reset.reset_n
		output wire         done,                    //    return.valid
		input  wire         stall                    //          .stall
	);

	cnn_top_internal cnn_top_internal_inst (
		.clock                   (clock),                   //     clock.clk
		.resetn                  (resetn),                  //     reset.reset_n
		.start                   (start),                   //      call.valid
		.busy                    (busy),                    //          .stall
		.done                    (done),                    //    return.valid
		.stall                   (stall),                   //          .stall
		.ddr_in1                 (ddr_in1),                 //   ddr_in1.data
		.ddr_w1                  (ddr_w1),                  //    ddr_w1.data
		.ddr_out1                (ddr_out1),                //  ddr_out1.data
		.param                   (param),                   //     param.data
		.ddr_scale               (ddr_scale),               // ddr_scale.data
		.avmm_1_rw_address       (avmm_1_rw_address),       // avmm_1_rw.address
		.avmm_1_rw_byteenable    (avmm_1_rw_byteenable),    //          .byteenable
		.avmm_1_rw_readdatavalid (avmm_1_rw_readdatavalid), //          .readdatavalid
		.avmm_1_rw_read          (avmm_1_rw_read),          //          .read
		.avmm_1_rw_readdata      (avmm_1_rw_readdata),      //          .readdata
		.avmm_1_rw_write         (avmm_1_rw_write),         //          .write
		.avmm_1_rw_writedata     (avmm_1_rw_writedata),     //          .writedata
		.avmm_1_rw_waitrequest   (avmm_1_rw_waitrequest),   //          .waitrequest
		.avmm_1_rw_burstcount    (avmm_1_rw_burstcount),    //          .burstcount
		.avmm_2_rw_address       (avmm_2_rw_address),       // avmm_2_rw.address
		.avmm_2_rw_byteenable    (avmm_2_rw_byteenable),    //          .byteenable
		.avmm_2_rw_readdatavalid (avmm_2_rw_readdatavalid), //          .readdatavalid
		.avmm_2_rw_read          (avmm_2_rw_read),          //          .read
		.avmm_2_rw_readdata      (avmm_2_rw_readdata),      //          .readdata
		.avmm_2_rw_write         (avmm_2_rw_write),         //          .write
		.avmm_2_rw_writedata     (avmm_2_rw_writedata),     //          .writedata
		.avmm_2_rw_waitrequest   (avmm_2_rw_waitrequest),   //          .waitrequest
		.avmm_2_rw_burstcount    (avmm_2_rw_burstcount),    //          .burstcount
		.avmm_3_rw_address       (avmm_3_rw_address),       // avmm_3_rw.address
		.avmm_3_rw_byteenable    (avmm_3_rw_byteenable),    //          .byteenable
		.avmm_3_rw_readdatavalid (avmm_3_rw_readdatavalid), //          .readdatavalid
		.avmm_3_rw_read          (avmm_3_rw_read),          //          .read
		.avmm_3_rw_readdata      (avmm_3_rw_readdata),      //          .readdata
		.avmm_3_rw_write         (avmm_3_rw_write),         //          .write
		.avmm_3_rw_writedata     (avmm_3_rw_writedata),     //          .writedata
		.avmm_3_rw_waitrequest   (avmm_3_rw_waitrequest),   //          .waitrequest
		.avmm_3_rw_burstcount    (avmm_3_rw_burstcount),    //          .burstcount
		.avmm_4_rw_address       (avmm_4_rw_address),       // avmm_4_rw.address
		.avmm_4_rw_byteenable    (avmm_4_rw_byteenable),    //          .byteenable
		.avmm_4_rw_readdatavalid (avmm_4_rw_readdatavalid), //          .readdatavalid
		.avmm_4_rw_read          (avmm_4_rw_read),          //          .read
		.avmm_4_rw_readdata      (avmm_4_rw_readdata),      //          .readdata
		.avmm_4_rw_write         (avmm_4_rw_write),         //          .write
		.avmm_4_rw_writedata     (avmm_4_rw_writedata),     //          .writedata
		.avmm_4_rw_waitrequest   (avmm_4_rw_waitrequest),   //          .waitrequest
		.avmm_4_rw_burstcount    (avmm_4_rw_burstcount),    //          .burstcount
		.avmm_5_rw_address       (avmm_5_rw_address),       // avmm_5_rw.address
		.avmm_5_rw_byteenable    (avmm_5_rw_byteenable),    //          .byteenable
		.avmm_5_rw_readdatavalid (avmm_5_rw_readdatavalid), //          .readdatavalid
		.avmm_5_rw_read          (avmm_5_rw_read),          //          .read
		.avmm_5_rw_readdata      (avmm_5_rw_readdata),      //          .readdata
		.avmm_5_rw_write         (avmm_5_rw_write),         //          .write
		.avmm_5_rw_writedata     (avmm_5_rw_writedata),     //          .writedata
		.avmm_5_rw_waitrequest   (avmm_5_rw_waitrequest),   //          .waitrequest
		.avmm_5_rw_burstcount    (avmm_5_rw_burstcount)     //          .burstcount
	);

endmodule
