// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// $Revision: #1 $
// $Date: 2018/07/18 $
// $Author: psgswbuild $

// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_arriagx_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

// ============================================================
// File Name: altera_streaming_sld_hub_controller_arriaiigx_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Arria II GX" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_arriaiigx_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	arriaii_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "arriaii_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_arriaiigx_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_arriaiigx_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_arriaiigx_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_arriaiigx_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigx_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigx_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigx_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigx_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigx_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigx_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_arriaiigz_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Arria II GZ" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_arriaiigz_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	arriaiigz_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "arriaiigz_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_arriaiigz_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_arriaiigz_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_arriaiigz_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_arriaiigz_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GZ"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GZ"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigz_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigz_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigz_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigz_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigz_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriaiigz_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_arriav_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Arria V" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = arriav_clkena 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_arriav_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	arriav_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk));
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "arriav_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_arriav_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_arriav_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_arriav_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_arriav_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria V"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriav_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriav_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriav_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriav_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriav_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_arriav_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_cycloneii_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// ============================================================
// File Name: altera_streaming_sld_hub_controller_cycloneiii_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Cyclone III" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" clkselect ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_cycloneiii_altclkctrl_altclkctrl
	( 
	clkselect,
	ena,
	inclk,
	outclk) ;
	input   [1:0]  clkselect;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0   [1:0]  clkselect;
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_clkctrl1_outclk;
	wire  [1:0]  clkselect_wire;
	wire  [3:0]  inclk_wire;

	cycloneiii_clkctrl   clkctrl1
	( 
	.clkselect(clkselect_wire),
	.ena(ena),
	.inclk(inclk_wire),
	.outclk(wire_clkctrl1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		clkctrl1.clock_type = "Global Clock",
		clkctrl1.ena_register_mode = "falling edge",
		clkctrl1.lpm_type = "cycloneiii_clkctrl";
	assign
		clkselect_wire = {clkselect},
		inclk_wire = {inclk},
		outclk = wire_clkctrl1_outclk;
endmodule //altera_streaming_sld_hub_controller_cycloneiii_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_cycloneiii_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [1:0] sub_wire1 = 2'h0;
	wire [2:0] sub_wire4 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire2 = inclk;
	wire [3:0] sub_wire3 = {sub_wire4, sub_wire2};

	altera_streaming_sld_hub_controller_cycloneiii_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_cycloneiii_altclkctrl_altclkctrl_component (
				.clkselect (sub_wire1),
				.ena (ena),
				.inclk (sub_wire3),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @clkselect 0 0 2 0 GND 0 0 2 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiii_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiii_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiii_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiii_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiii_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiii_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Cyclone III LS" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" clkselect ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl_altclkctrl
	( 
	clkselect,
	ena,
	inclk,
	outclk) ;
	input   [1:0]  clkselect;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0   [1:0]  clkselect;
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_clkctrl1_outclk;
	wire  [1:0]  clkselect_wire;
	wire  [3:0]  inclk_wire;

	cycloneiiils_clkctrl   clkctrl1
	( 
	.clkselect(clkselect_wire),
	.ena(ena),
	.inclk(inclk_wire),
	.outclk(wire_clkctrl1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		clkctrl1.clock_type = "Global Clock",
		clkctrl1.ena_register_mode = "falling edge",
		clkctrl1.lpm_type = "cycloneiiils_clkctrl";
	assign
		clkselect_wire = {clkselect},
		inclk_wire = {inclk},
		outclk = wire_clkctrl1_outclk;
endmodule //altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [1:0] sub_wire1 = 2'h0;
	wire [2:0] sub_wire4 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire2 = inclk;
	wire [3:0] sub_wire3 = {sub_wire4, sub_wire2};

	altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl_altclkctrl_component (
				.clkselect (sub_wire1),
				.ena (ena),
				.inclk (sub_wire3),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III LS"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III LS"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @clkselect 0 0 2 0 GND 0 0 2 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneiiils_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_cycloneive_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Cyclone IV E" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" clkselect ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_cycloneive_altclkctrl_altclkctrl
	( 
	clkselect,
	ena,
	inclk,
	outclk) ;
	input   [1:0]  clkselect;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0   [1:0]  clkselect;
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_clkctrl1_outclk;
	wire  [1:0]  clkselect_wire;
	wire  [3:0]  inclk_wire;

	cycloneive_clkctrl   clkctrl1
	( 
	.clkselect(clkselect_wire),
	.ena(ena),
	.inclk(inclk_wire),
	.outclk(wire_clkctrl1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		clkctrl1.clock_type = "Global Clock",
		clkctrl1.ena_register_mode = "falling edge",
		clkctrl1.lpm_type = "cycloneive_clkctrl";
	assign
		clkselect_wire = {clkselect},
		inclk_wire = {inclk},
		outclk = wire_clkctrl1_outclk;
endmodule //altera_streaming_sld_hub_controller_cycloneive_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_cycloneive_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [1:0] sub_wire1 = 2'h0;
	wire [2:0] sub_wire4 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire2 = inclk;
	wire [3:0] sub_wire3 = {sub_wire4, sub_wire2};

	altera_streaming_sld_hub_controller_cycloneive_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_cycloneive_altclkctrl_altclkctrl_component (
				.clkselect (sub_wire1),
				.ena (ena),
				.inclk (sub_wire3),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @clkselect 0 0 2 0 GND 0 0 2 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneive_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneive_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneive_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneive_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneive_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneive_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Cyclone IV GX" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" clkselect ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl_altclkctrl
	( 
	clkselect,
	ena,
	inclk,
	outclk) ;
	input   [1:0]  clkselect;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0   [1:0]  clkselect;
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_clkctrl1_outclk;
	wire  [1:0]  clkselect_wire;
	wire  [3:0]  inclk_wire;

	cycloneiv_clkctrl   clkctrl1
	( 
	.clkselect(clkselect_wire),
	.ena(ena),
	.inclk(inclk_wire),
	.outclk(wire_clkctrl1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		clkctrl1.clock_type = "Global Clock",
		clkctrl1.ena_register_mode = "falling edge",
		clkctrl1.lpm_type = "cycloneiv_clkctrl";
	assign
		clkselect_wire = {clkselect},
		inclk_wire = {inclk},
		outclk = wire_clkctrl1_outclk;
endmodule //altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [1:0] sub_wire1 = 2'h0;
	wire [2:0] sub_wire4 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire2 = inclk;
	wire [3:0] sub_wire3 = {sub_wire4, sub_wire2};

	altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl_altclkctrl_component (
				.clkselect (sub_wire1),
				.ena (ena),
				.inclk (sub_wire3),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @clkselect 0 0 2 0 GND 0 0 2 0
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cycloneivgx_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_cyclonev_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Cyclone V" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = cyclonev_clkena 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_cyclonev_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	cyclonev_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk));
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "cyclonev_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_cyclonev_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_cyclonev_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_cyclonev_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_cyclonev_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cyclonev_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cyclonev_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cyclonev_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cyclonev_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cyclonev_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_cyclonev_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_stratixii_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// ============================================================
// File Name: altera_streaming_sld_hub_controller_stratixiii_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Stratix III" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_stratixiii_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	stratixiii_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "stratixiii_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_stratixiii_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_stratixiii_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_stratixiii_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_stratixiii_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiii_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiii_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiii_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiii_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiii_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiii_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_stratixiv_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Stratix IV" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = clkctrl 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_stratixiv_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	// wire [1:0]  clkselect;

	stratixiv_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk)
	// synopsys translate_off
	,
	.devclrn(1'b1),
	.devpor(1'b1)
	// synopsys translate_on
	);
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "stratixiv_clkena";
	assign
		// clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_stratixiv_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_stratixiv_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_stratixiv_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_stratixiv_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiv_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiv_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiv_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiv_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiv_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixiv_altclkctrl_bb.v FALSE
// megafunction wizard: %ALTCLKCTRL%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altclkctrl 

// ============================================================
// File Name: altera_streaming_sld_hub_controller_stratixv_altclkctrl.v
// Megafunction Name(s):
// 			altclkctrl
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.0 Internal Build 65 11/10/2011 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


//altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Stratix V" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 12.0 cbx_altclkbuf 2011:11:10:21:13:25:SJ cbx_cycloneii 2011:11:10:21:13:25:SJ cbx_lpm_add_sub 2011:11:10:21:13:25:SJ cbx_lpm_compare 2011:11:10:21:13:25:SJ cbx_lpm_decode 2011:11:10:21:13:25:SJ cbx_lpm_mux 2011:11:10:21:13:25:SJ cbx_mgl 2011:11:10:21:21:46:SJ cbx_stratix 2011:11:10:21:13:25:SJ cbx_stratixii 2011:11:10:21:13:25:SJ cbx_stratixiii 2011:11:10:21:13:25:SJ cbx_stratixv 2011:11:10:21:13:25:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463


//synthesis_resources = stratixv_clkena 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_stratixv_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) ;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	stratixv_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk));
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "stratixv_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //altera_streaming_sld_hub_controller_stratixv_altclkctrl_altclkctrl
//VALID FILE


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_streaming_sld_hub_controller_stratixv_altclkctrl (
	ena,
	inclk,
	outclk);

	input	  ena;
	input	  inclk;
	output	  outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  sub_wire0;
	wire [2:0] sub_wire3 = 3'h0;
	wire  outclk = sub_wire0;
	wire  sub_wire1 = inclk;
	wire [3:0] sub_wire2 = {sub_wire3, sub_wire1};

	altera_streaming_sld_hub_controller_stratixv_altclkctrl_altclkctrl	altera_streaming_sld_hub_controller_stratixv_altclkctrl_altclkctrl_component (
				.ena (ena),
				.inclk (sub_wire2),
				.outclk (sub_wire0));

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: clock_inputs NUMERIC "1"
// Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "OFF"
// Retrieval info: CONSTANT: clock_type STRING "Global Clock"
// Retrieval info: USED_PORT: ena 0 0 0 0 INPUT VCC "ena"
// Retrieval info: USED_PORT: inclk 0 0 0 0 INPUT NODEFVAL "inclk"
// Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
// Retrieval info: CONNECT: @ena 0 0 0 0 ena 0 0 0 0
// Retrieval info: CONNECT: @inclk 0 0 3 1 GND 0 0 3 0
// Retrieval info: CONNECT: @inclk 0 0 1 0 inclk 0 0 0 0
// Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixv_altclkctrl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixv_altclkctrl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixv_altclkctrl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixv_altclkctrl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixv_altclkctrl_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_streaming_sld_hub_controller_stratixv_altclkctrl_bb.v FALSE

//altclkctrl CBX_SINGLE_OUTPUT_FILE="ON" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Arria 10" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="OFF" ena inclk outclk
//VERSION_BEGIN 15.1 cbx_altclkbuf 2015:10:14:18:59:15:SJ cbx_cycloneii 2015:10:14:18:59:15:SJ cbx_lpm_add_sub 2015:10:14:18:59:15:SJ cbx_lpm_compare 2015:10:14:18:59:15:SJ cbx_lpm_decode 2015:10:14:18:59:15:SJ cbx_lpm_mux 2015:10:14:18:59:15:SJ cbx_mgl 2015:10:21:19:02:34:SJ cbx_nadder 2015:10:14:18:59:15:SJ cbx_stratix 2015:10:14:18:59:15:SJ cbx_stratixii 2015:10:14:18:59:15:SJ cbx_stratixiii 2015:10:14:18:59:15:SJ cbx_stratixv 2015:10:14:18:59:15:SJ  VERSION_END
// synthesis VERILOG_INPUT_VERSION VERILOG_2001
// altera message_off 10463



// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
//  Your use of Altera Corporation's design tools, logic functions 
//  and other software and tools, and its AMPP partner logic 
//  functions, and any output files from any of the foregoing 
//  (including device programming or simulation files), and any 
//  associated documentation or information are expressly subject 
//  to the terms and conditions of the Altera Program License 
//  Subscription Agreement, the Altera Quartus Prime License Agreement,
//  the Altera MegaCore Function License Agreement, or other 
//  applicable license agreement, including, without limitation, 
//  that your use is for the sole purpose of programming logic 
//  devices manufactured by Altera and sold by Altera or its 
//  authorized distributors.  Please refer to the applicable 
//  agreement for further details.



//synthesis_resources = twentynm_clkena 1 
//synopsys translate_off
`timescale 1 ps / 1 ps
//synopsys translate_on
module  altera_streaming_sld_hub_controller_arria10_altclkctrl_altclkctrl
	( 
	ena,
	inclk,
	outclk) /* synthesis synthesis_clearbox=1 */;
	input   ena;
	input   [3:0]  inclk;
	output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1   ena;
	tri0   [3:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire  wire_sd1_outclk;
	wire [1:0]  clkselect;

	twentynm_clkena   sd1
	( 
	.ena(ena),
	.enaout(),
	.inclk(inclk[0]),
	.outclk(wire_sd1_outclk));
	defparam
		sd1.clock_type = "Global Clock",
		sd1.ena_register_mode = "falling edge",
		sd1.lpm_type = "twentynm_clkena";
	assign
		clkselect = {2{1'b0}},
		outclk = wire_sd1_outclk;
endmodule //a10_altclk_altclkctrl_151_6g5aioa_sub
//VALID FILE // (C) 2001-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.



// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module  altera_streaming_sld_hub_controller_arria10_altclkctrl  (
    ena,
    inclk,
    outclk);

    input    ena;
    input    inclk;
    output   outclk;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
    tri1     ena;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

    wire  sub_wire0;
    wire  outclk;
    wire  sub_wire1;
    wire [3:0] sub_wire2;
    wire [2:0] sub_wire3;

    assign  outclk = sub_wire0;
    assign  sub_wire1 = inclk;
    assign sub_wire2[3:0] = {sub_wire3, sub_wire1};
    assign sub_wire3[2:0] = 3'h0;

    altera_streaming_sld_hub_controller_arria10_altclkctrl_altclkctrl  altera_streaming_sld_hub_controller_arria10_altclkctrl_altclkctrl_component (
                .ena (ena),
                .inclk (sub_wire2),
                .outclk (sub_wire0));

endmodule
